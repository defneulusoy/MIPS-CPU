//Property of Prof. J. Marpaung and Northeastern University
//Not to be distributed elsewhere without a written consent from Prof. J. Marpaung
//All Rights Reserved
`timescale 1ns/10ps
module cpu5_testbench();
reg [31:0] instrbus;
reg [31:0] instrbusin[0:99];
wire [31:0] iaddrbus, daddrbus;
reg [31:0] iaddrbusout[0:99], daddrbusout[0:99];
wire [31:0] databus;
  reg [31:0] databusk, databusin[0:99], databusout[0:99];
reg clk, reset;
reg clkd;
reg [31:0] dontcare;
reg [24*8:1] iname[0:99];
integer error, k, ntests;
parameter Rformat = 6'b000000;
parameter ADDI = 6'b000011;
parameter SUBI = 6'b000010;
parameter XORI = 6'b000001;
parameter ANDI = 6'b001111;
parameter ORI = 6'b001100;
parameter LW = 6'b011110;
parameter SW = 6'b011111;
parameter BEQ = 6'b110000;
parameter BNE = 6'b110001;
parameter ADD = 6'b000011;
parameter SUB = 6'b000010;
parameter XOR = 6'b000001;
parameter AND = 6'b000111;
parameter OR = 6'b000100;
parameter SLT = 6'b110110;
parameter SLE = 6'b110111;
cpu5
dut(.reset(reset),.clk(clk),.iaddrbus(iaddrbus),.ibus(instrbus),.daddrbus(daddrbus),.databus(databus));
initial begin
// This test file runs the following program.
iname[0] = "ADDI R20, R0, #-1";
iname[1] = "ADDI R21, R0, #1";
iname[2] = "ADDI R22, R0, #2";
iname[3] = "LW R24, 0(R20)";
iname[4] = "LW R25, 0(R21)";
iname[5] = "SW 1000(R22), R20";
iname[6] = "SW 2(R0), R21";
iname[7] = "ADD R26, R24, R25";
iname[8] = "SUBI R17, R24, 6420";
iname[9] = "SUB R27, R24, R25";
iname[10] = "ANDI R18, R24, #0";
iname[11] = "AND R28, R24, R0";
iname[12] = "XORI R19, R24, 6420";
iname[13] = "XOR R29, R24, R25";
iname[14] = "ORI R20, R24, 6420";
iname[15] = "OR R30, R24, R25";
iname[16] = "SW 0(R26), R26";
iname[17] = "SW 0(R17), R27";
iname[18] = "SW 1000(R18), R28";
iname[19] = "SW 0(R19), R29";
iname[20] = "SW 0(R20), R30";
iname[21] = "SLT R1, R0, R21"; // Setting R1 to 32'h00000001 (since, R0 < R21).
iname[22] = "ADDI R5, R0, #1";
iname[23] = "ADDI R6, R0, #1";
  iname[24] = "BNE R0, R1, #10"; // Branching to (32'h00000060 + 32'h00000004 + 32'h00000028 = 32'h0000008C) since, R0 != R1.
iname[25] = "ADDI R8, R0, #1"; // Delay Slot
//Branched Location - 32'h0000008C //
iname[26] = "SLE R2, R0, R0"; // Setting R2 to 32'h00000001 (since, R0 = R0).
iname[27] = "NOP";
iname[28] = "NOP";
iname[29] = "BEQ R0, R2, #25"; // NOT Branching since, R2 != R0.
iname[30] = "NOP"; // Delay Slot
  iname[31] = "BEQ R2, R2, #10"; // Branching to (32h'0000000A0 + 32'h00000004 + 32'h00000028 = 32'h000000CC)
iname[32] = "ADDI R20, R0, #1"; // Delay Slot
//Branched Location - 32'h000000CC //
iname[33] = "NOP";
iname[34] = "NOP";
iname[35] = "NOP";
  
iname[36] = "ORI R20, R0, #-2";
iname[37] = "XORI R21, R0, #2";
iname[38] = "XORI R22, R0, #4";
iname[39] = "LW R24, 0(R20)";
iname[40] = "LW R25, 0(R21)";
iname[41] = "SW 1000(R22), R20";
iname[42] = "SW 2(R0), R21";
iname[43] = "SUB R26, R24, R25";
iname[44] = "SUBI R17, R24, 1010";
iname[45] = "ADD R27, R24, R25";
iname[46] = "ORI R18, R24, #0";
iname[47] = "XOR R28, R24, R0";
iname[48] = "ADDI R19, R24, F0F0";
iname[49] = "ADD R29, R24, R25";
iname[50] = "ADDI R20, R24, AAAA";
iname[51] = "XOR R30, R24, R25";
iname[52] = "SW 0(R26), R26";
iname[53] = "SW 0(R17), R27";
iname[54] = "SW 1000(R18), R28";
iname[55] = "SW 0(R19), R29";
iname[56] = "SW 0(R20), R30";
iname[57] = "SLE R1, R0, R21";      
iname[58] = "ORI R5, R0, #4";
iname[59] = "SUBI R6, R0, #2";
iname[60] = "BNE R0, R1, #20";
iname[61] = "XORI R8, R0, #00FF";
iname[62] = "SLT R2, R0, R0";
iname[63] = "NOP";
iname[64] = "NOP";
iname[65] = "BEQ R0, R2, #10";
iname[66] = "NOP";
iname[67] = "BEQ R2, R2, #80";
iname[68] = "ORI R20, R0, #4444";
iname[69] = "";
iname[70] = "";
iname[71] = "";
iname[72] = "";
iname[73] = "";
iname[74] = "";
iname[75] = "";
iname[76] = "";
iname[77] = "";
iname[78] = "";
iname[79] = "";
iname[80] = "";
iname[81] = "";
iname[82] = "";
iname[83] = "";
iname[84] = "";
iname[85] = "";
iname[86] = "";
iname[87] = "";
iname[88] = "";
iname[89] = "";
iname[90] = "";
iname[91] = "";
iname[92] = "";
iname[93] = "";
iname[94] = "";
iname[95] = "";
iname[96] = "";
iname[97] = "";
iname[98] = "";
iname[99] = "";

  
dontcare = 32'hx;
//* ADDI R20, R0, #-1
iaddrbusout[0] = 32'h00000000;
// opcode source1 dest Immediate...
instrbusin[0]={ADDI, 5'b00000, 5'b10100, 16'hFFFF};
daddrbusout[0] = dontcare;
databusin[0] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[0] = dontcare;
//* ADDI R21, R0, #1
iaddrbusout[1] = 32'h00000004;
// opcode source1 dest Immediate...
instrbusin[1]={ADDI, 5'b00000, 5'b10101, 16'h0001};
daddrbusout[1] = dontcare;
databusin[1] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[1] = dontcare;
//* ADDI R22, R0, #2
iaddrbusout[2] = 32'h00000008;
// opcode source1 dest Immediate...
instrbusin[2]={ADDI, 5'b00000, 5'b10110, 16'h0002};
daddrbusout[2] = dontcare;
databusin[2] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[2] = dontcare;
//* LW R24, 0(R20)
iaddrbusout[3] = 32'h0000000C;
// opcode source1 dest Immediate...
instrbusin[3]={LW, 5'b10100, 5'b11000, 16'h0000};
daddrbusout[3] = 32'hFFFFFFFF;
databusin[3] = 32'hCCCCCCCC;
databusout[3] = dontcare;
//* LW R25, 0(R21)
iaddrbusout[4] = 32'h00000010;
// opcode source1 dest Immediate...
instrbusin[4]={LW, 5'b10101, 5'b11001, 16'h0000};
daddrbusout[4] = 32'h00000001;
databusin[4] = 32'hAAAAAAAA;
databusout[4] = dontcare;
//* SW 1000(R22), R20
iaddrbusout[5] = 32'h00000014;
// opcode source1 dest Immediate...
instrbusin[5]={SW, 5'b10110, 5'b10100, 16'h1000};
daddrbusout[5] = 32'h00001002;
databusin[5] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[5] = 32'hFFFFFFFF;
//* SW 2(R0), R21
iaddrbusout[6] = 32'h00000018;
// opcode source1 dest Immediate...
instrbusin[6]={SW, 5'b00000, 5'b10101, 16'h0002};
daddrbusout[6] = 32'h00000002;
databusin[6] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[6] = 32'h00000001;
//* ADD R26, R24, R25
iaddrbusout[7] = 32'h0000001C;
// opcode source1 source2 dest shift Function...
instrbusin[7]={Rformat, 5'b11000, 5'b11001, 5'b11010, 5'b00000, ADD};
daddrbusout[7] = dontcare;
databusin[7] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[7] = dontcare;
//* SUBI R17, R24, 6420
iaddrbusout[8] = 32'h00000020;
// opcode source1 dest Immediate...
instrbusin[8]={SUBI, 5'b11000, 5'b10001, 16'h6420};
daddrbusout[8] = dontcare;
databusin[8] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[8] = dontcare;
//* SUB R27, R24, R25
iaddrbusout[9] = 32'h00000024;
// opcode source1 source2 dest shift Function...
instrbusin[9]={Rformat, 5'b11000, 5'b11001, 5'b11011, 5'b00000, SUB};
daddrbusout[9] = dontcare;
databusin[9] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[9] = dontcare;
//* ANDI R18, R24, #0
iaddrbusout[10] = 32'h00000028;
// opcode source1 dest Immediate...
instrbusin[10]={ANDI, 5'b11000, 5'b10010, 16'h0000};
daddrbusout[10] = dontcare;
databusin[10] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[10] = dontcare;
//* AND R28, R24, R0
iaddrbusout[11] = 32'h0000002C;
// opcode source1 source2 dest shift Function...
instrbusin[11]={Rformat, 5'b11000, 5'b00000, 5'b11100, 5'b00000, AND};
daddrbusout[11] = dontcare;
databusin[11] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[11] = dontcare;
//* XORI R19, R24, 6420
iaddrbusout[12] = 32'h00000030;
// opcode source1 dest Immediate...
instrbusin[12]={XORI, 5'b11000, 5'b10011, 16'h6420};
daddrbusout[12] = dontcare;
databusin[12] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[12] = dontcare;
//* XOR R29, R24, R25
iaddrbusout[13] = 32'h00000034;
// opcode source1 source2 dest shift Function...
instrbusin[13]={Rformat, 5'b11000, 5'b11001, 5'b11101, 5'b00000, XOR};
daddrbusout[13] = dontcare;
databusin[13] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[13] = dontcare;
//* ORI R20, R24, 6420
iaddrbusout[14] = 32'h00000038;
// opcode source1 dest Immediate...
instrbusin[14]={ORI, 5'b11000, 5'b10100, 16'h6420};
daddrbusout[14] = dontcare;
databusin[14] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[14] = dontcare;
//* OR R30, R24, R25
iaddrbusout[15] = 32'h0000003C;
// opcode source1 source2 dest shift Function...
instrbusin[15]={Rformat, 5'b11000, 5'b11001, 5'b11110, 5'b00000, OR};
daddrbusout[15] = dontcare;
databusin[15] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[15] = dontcare;
//* SW 0(R26), R26
iaddrbusout[16] = 32'h00000040;
// opcode source1 dest Immediate...
instrbusin[16]={SW, 5'b11010, 5'b11010, 16'h0000};
daddrbusout[16] = 32'h77777776;
databusin[16] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[16] = 32'h77777776;
//18* SW 0(R17), R27
iaddrbusout[17] = 32'h00000044;
// opcode source1 dest Immediate...
instrbusin[17]={SW, 5'b10001, 5'b11011, 16'h0000};
daddrbusout[17] = 32'hCCCC68AC;
databusin[17] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[17] = 32'h22222222;
//19* SW 1000(R18), R28
iaddrbusout[18] = 32'h00000048;
// opcode source1 dest Immediate...
instrbusin[18]={SW, 5'b10010, 5'b11100, 16'h1000};
daddrbusout[18] = 32'h00001000;
databusin[18] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[18] = 32'h00000000;
//20* SW 0(R19), R29
iaddrbusout[19] = 32'h0000004C;
// opcode source1 dest Immediate...
instrbusin[19]={SW, 5'b10011, 5'b11101, 16'h0000};
daddrbusout[19] = 32'hCCCCA8EC;
databusin[19] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[19] = 32'h66666666;
//21* SW 0(R20), R30
iaddrbusout[20] = 32'h00000050;
// opcode source1 dest Immediate...
instrbusin[20]={SW, 5'b10100, 5'b11110, 16'h0000};
daddrbusout[20] = 32'hCCCCECEC;
databusin[20] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[20] = 32'hEEEEEEEE;
//22* SLT R1, R0, R21
iaddrbusout[21] = 32'h00000054;
// opcode source1 source2 dest shift Function...
instrbusin[21]={Rformat, 5'b00000, 5'b10101, 5'b00001, 5'b00000, SLT};
daddrbusout[21] = dontcare;
databusin[21] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[21] = dontcare;
//* ADDI R5, R0, #1
iaddrbusout[22] = 32'h00000058;
// opcode source1 dest Immediate...
instrbusin[22]={ADDI, 5'b00000, 5'b00101, 16'h0001};
daddrbusout[22] = dontcare;
databusin[22] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[22] = dontcare;
//* ADDI R6, R0, #1
iaddrbusout[23] = 32'h0000005C;
// opcode source1 dest Immediate...
instrbusin[23]={ADDI, 5'b00000, 5'b00110, 16'h0001};
daddrbusout[23] = dontcare;
databusin[23] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[23] = dontcare;
//* BNE R0, R1, #10
iaddrbusout[24] = 32'h00000060;
// opcode source1 dest Immediate...
instrbusin[24]={BNE, 5'b00001, 5'b00000, 16'h000A};
daddrbusout[24] = dontcare;
databusin[24] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[24] = dontcare;
//* ADDI R8, R0, #1
iaddrbusout[25] = 32'h00000064;
// opcode source1 dest Immediate...
instrbusin[25]={ADDI, 5'b00000, 5'b01000, 16'h0001};
daddrbusout[25] = dontcare;
databusin[25] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[25] = dontcare;
//* SLE R2, R0, R0
iaddrbusout[26] = 32'h0000008C;
// opcode source1 source2 dest shift Function...
instrbusin[26]={Rformat, 5'b00000, 5'b00000, 5'b00010, 5'b00000, SLE};
daddrbusout[26] = dontcare;
databusin[26] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[26] = dontcare;
//* NOP
iaddrbusout[27] = 32'h00000090;
// oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[27] = 32'b00000000000000000000000000000000;
daddrbusout[27] = dontcare;
databusin[27] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[27] = dontcare;
//* NOP
iaddrbusout[28] = 32'h00000094;
// oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[28] = 32'b00000000000000000000000000000000;
daddrbusout[28] = dontcare;
databusin[28] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[28] = dontcare;
//* BEQ R0, R2, #25
iaddrbusout[29] = 32'h00000098;
// opcode source1 dest Immediate...
instrbusin[29]={BEQ, 5'b00010, 5'b00000, 16'h0019};
daddrbusout[29] = dontcare;
databusin[29] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[29] = dontcare;
//* NOP
iaddrbusout[30] = 32'h0000009C;
// oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[30] = 32'b00000000000000000000000000000000;
daddrbusout[30] = dontcare;
databusin[30] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[30] = dontcare;
//* BEQ R2, R2, #10
iaddrbusout[31] = 32'h000000A0;
// opcode source1 dest Immediate...
instrbusin[31]={BEQ, 5'b00010, 5'b00010, 16'h000A};
daddrbusout[31] = dontcare;
databusin[31] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[31] = dontcare;
//* ADDI R20, R0, #1
iaddrbusout[32] = 32'h000000A4;
// opcode source1 dest Immediate...
instrbusin[32]={ADDI, 5'b00000, 5'b10100, 16'h0001};
daddrbusout[32] = dontcare;
databusin[32] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[32] = dontcare;
//* NOP
iaddrbusout[33] = 32'h000000CC;
// oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[33] = 32'b00000000000000000000000000000000;
daddrbusout[33] = dontcare;
databusin[33] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[33] = dontcare;
//* NOP
iaddrbusout[34] = 32'h000000D0;
// oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[34] = 32'b00000000000000000000000000000000;
daddrbusout[34] = dontcare;
databusin[34] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[34] = dontcare;
//* NOP
iaddrbusout[35] = 32'h000000D4;
// oooooosssssdddddiiiiiiiiiiiiiiii
instrbusin[35] = 32'b00000000000000000000000000000000;
daddrbusout[35] = dontcare;
databusin[35] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[35] = dontcare;
  
  
//* ORI R20, R0, #-2
iaddrbusout[36] = 32'b00000000000000000000000011011000;
instrbusin[36]={ORI, 5'b00000, 5'b10100, 16'hFFFE};
daddrbusout[36] = dontcare;
databusin[36] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[36] = dontcare;
  
//* XORI R21, R0, #2
iaddrbusout[37] = 32'b0000000000000000000000011011100;
instrbusin[37]={XORI, 5'b00000, 5'b10101, 16'h0002};
daddrbusout[37] = dontcare;
databusin[37] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[37] = dontcare;
  
//* XORI R22, R0, #4
iaddrbusout[38] = 32'b00000000000000000000000011100000;
instrbusin[38]={XORI, 5'b00000, 5'b10110, 16'h0004};
daddrbusout[38] = dontcare;
databusin[38] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[38] = dontcare;
  
//* LW R24, 0(R20), R24 = -2
iaddrbusout[39] = 32'b00000000000000000000000011100100;
instrbusin[39]={LW, 5'b10100, 5'b11000, 16'h0000};
daddrbusout[39] = 32'hFFFFFFFE;
databusin[39] = 32'hCCCCCCCC;
databusout[39] = dontcare;
  
//* LW R25, 0(R21) R25 = 2
iaddrbusout[40] = 32'b 00000000000000000000000011101000;
instrbusin[40]={LW, 5'b10101, 5'b11001, 16'h0000};
daddrbusout[40] = 32'h00000002;
databusin[40] = 32'hAAAAAAAA;
databusout[40] = dontcare;
  
//* SW 1000(R22), R20
iaddrbusout[41] = 32'b 00000000000000000000000011101100;
instrbusin[41]={SW, 5'b10110, 5'b10100, 16'h1000};
daddrbusout[41] = 32'h00001004;
databusin[41] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[41] = 32'hFFFFFFFE;
  
//* SW 2(R0), R21
iaddrbusout[42] = 32'b00000000000000000000000011110000;
instrbusin[42]={SW, 5'b00000, 5'b10101, 16'h0002};
daddrbusout[42] = 32'h00000002;
databusin[42] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[42] = 32'h00000002;
  
//* SUB R26, R24, R25
iaddrbusout[43] = 32'b00000000000000000000000011110100;
instrbusin[43]={Rformat, 5'b11000, 5'b11001, 5'b11010, 5'b00000, SUB};
daddrbusout[43] = dontcare;
databusin[43] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[43] = dontcare;
  
//* SUBI R17, R24, 1010
iaddrbusout[44] = 32'b00000000000000000000000011111000;
instrbusin[44]={SUBI, 5'b11000, 5'b10001, 16'h1010};
daddrbusout[44] = dontcare;
databusin[44] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[44] = dontcare;
  
//* ADD R27, R24, R25
iaddrbusout[45] = 32'b00000000000000000000000011111100;
instrbusin[45]={Rformat, 5'b11000, 5'b11001, 5'b11011, 5'b00000, ADD};
daddrbusout[45] = dontcare;
databusin[45] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[45] = dontcare;
  
//* ORI R18, R24, #0
iaddrbusout[46] = 32'b00000000000000000000000100000000;
instrbusin[46]={ORI, 5'b11000, 5'b10010, 16'h0000};
daddrbusout[46] = dontcare;
databusin[46] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[46] = dontcare;
  
//* XOR R28, R24, R0
iaddrbusout[47] = 32'b00000000000000000000000100000100;
instrbusin[47]={Rformat, 5'b11000, 5'b00000, 5'b11100, 5'b00000, XOR};
daddrbusout[47] = dontcare;
databusin[47] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[47] = dontcare;
  
//* ADDI R19, R24, F0F0
iaddrbusout[48] = 32'b00000000000000000000000100001000;
instrbusin[48]={ADDI, 5'b11000, 5'b10011, 16'hF0F0};
daddrbusout[48] = dontcare;
databusin[48] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[48] = dontcare;
  
//* ADD R29, R24, R25
iaddrbusout[49] = 32'b00000000000000000000000100001100;
instrbusin[49]={Rformat, 5'b11000, 5'b11001, 5'b11101, 5'b00000, ADD};
daddrbusout[49] = dontcare;
databusin[49] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[49] = dontcare;
  
//* ADDI R20, R24, AAAA
iaddrbusout[50] = 32'b00000000000000000000000100010000;
instrbusin[50]={ADDI, 5'b11000, 5'b10100, 16'hAAAA};
daddrbusout[50] = dontcare;
databusin[50] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[50] = dontcare;
  
//* XOR R30, R24, R25
iaddrbusout[51] = 32'b00000000000000000000000100010100;
instrbusin[51]={Rformat, 5'b11000, 5'b11001, 5'b11110, 5'b00000, XOR};
daddrbusout[51] = dontcare;
databusin[51] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[51] = dontcare;
  
//* SW 0(R26), R26
iaddrbusout[52] = 32'b00000000000000000000000100011000;
instrbusin[52]={SW, 5'b11010, 5'b11010, 16'h0000};
daddrbusout[52] = 32'b00100010001000100010001000100010;
databusin[52] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[52] = 32'b00100010001000100010001000100010;
  
//18* SW 0(R17), R27
iaddrbusout[53] = 32'b00000000000000000000000100011100;
instrbusin[53]={SW, 5'b10001, 5'b11011, 16'h0000};
daddrbusout[53] = 32'b11001100110011001011110010111100;
databusin[53] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[53] = 32'b01110111011101110111011101110110;
  
//19* SW 1000(R18), R28
iaddrbusout[54] = 32'b00000000000000000000000100100000;
instrbusin[54]={SW, 5'b10010, 5'b11100, 16'h1000};
daddrbusout[54] = 32'b11001100110011001101110011001100;
databusin[54] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[54] = 32'b11001100110011001100110011001100;
  
//20* SW 0(R19), R29
iaddrbusout[55] = 32'b00000000000000000000000100100100;
instrbusin[55]={SW, 5'b10011, 5'b11101, 16'h0000};
daddrbusout[55] = 32'b11001100110011001011110110111100;
databusin[55] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[55] = 32'b01110111011101110111011101110110;
  
//21* SW 0(R20), R30
iaddrbusout[56] = 32'b00000000000000000000000100101000;
instrbusin[56]={SW, 5'b10100, 5'b11110, 16'h0000};
daddrbusout[56] = 32'b11001100110011000111011101110110;
databusin[56] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[56] = 32'b01100110011001100110011001100110;
  
//22* SLE R1, R0, R21
iaddrbusout[57] = 32'b00000000000000000000000100101100;
instrbusin[57]={Rformat, 5'b00000, 5'b10101, 5'b00001, 5'b00000, SLE};
daddrbusout[57] = dontcare;
databusin[57] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[57] = dontcare;
  
//* ORI R5, R0, #4
iaddrbusout[58] = 32'b00000000000000000000000100110000;
instrbusin[58]={ORI, 5'b00000, 5'b00101, 16'h0004};
daddrbusout[58] = dontcare;
databusin[58] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[58] = dontcare;
  
//* SUBI R6, R0, #2
iaddrbusout[59] = 32'b00000000000000000000000100110100;
instrbusin[59]={SUBI, 5'b00000, 5'b00110, 16'h0002};
daddrbusout[59] = dontcare;
databusin[59] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[59] = dontcare;
  
//* BNE R0, R1, #20
iaddrbusout[60] = 32'b00000000000000000000000100111000;
instrbusin[60]={BNE, 5'b00001, 5'b00000, 16'h0014};
daddrbusout[60] = dontcare;
databusin[60] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[60] = dontcare;
  
//* XORI R8, R0, #00FF
iaddrbusout[61] = 32'b00000000000000000000000100111100;
instrbusin[61]={XORI, 5'b00000, 5'b01000, 16'h00FF};
daddrbusout[61] = dontcare;
databusin[61] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[61] = dontcare;
  
//* SLT R2, R0, R0
iaddrbusout[62] = 32'b00000000000000000000000110001100;
instrbusin[62]={Rformat, 5'b00000, 5'b00000, 5'b00010, 5'b00000, SLT};
daddrbusout[62] = dontcare;
databusin[62] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[62] = dontcare;
  
//* NOP
iaddrbusout[63] = 32'b00000000000000000000000110010000;
instrbusin[63] = 32'b00000000000000000000000000000000;
daddrbusout[63] = dontcare;
databusin[63] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[63] = dontcare;
  
//* NOP
iaddrbusout[64] = 32'b00000000000000000000000110010100;
instrbusin[64] = 32'b00000000000000000000000000000000;
daddrbusout[64] = dontcare;
databusin[64] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[64] = dontcare;
  
//* BEQ R0, R2, #10
iaddrbusout[65] = 32'b00000000000000000000000110011000;
instrbusin[65]={BEQ, 5'b00010, 5'b00000, 16'h000A};
daddrbusout[65] = dontcare;
databusin[65] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[65] = dontcare;
  
//* NOP
iaddrbusout[66] = 32'b00000000000000000000000110011100;
instrbusin[66] = 32'b00000000000000000000000000000000;
daddrbusout[66] = dontcare;
databusin[66] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[66] = dontcare;
  
//* BEQ R2, R2, #80
iaddrbusout[67] = 32'b00000000000000000000000111000100;
instrbusin[67]={BEQ, 5'b00010, 5'b00010, 16'h0050};
daddrbusout[67] = dontcare;
databusin[67] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[67] = dontcare;
  
//* ORI R20, R0, #4444
iaddrbusout[68] = 32'b00000000000000000000000111001000;
instrbusin[68]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[68] = dontcare;
databusin[68] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[68] = dontcare;

iaddrbusout[69] = 32'b00000000000000000000001100001000;
instrbusin[69]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[69] = dontcare;
databusin[69] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[69] = dontcare;  

iaddrbusout[70] = 32'b00000000000000000000001100001100;
instrbusin[70]={SUBI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[70] = dontcare;
databusin[70] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[70] = dontcare;

iaddrbusout[71] = 32'b00000000000000000000001100010000;
instrbusin[71]={ORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[71] = dontcare;
databusin[71] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[71] = dontcare;

iaddrbusout[72] = 32'b00000000000000000000001100010100;
instrbusin[72]={XORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[72] = dontcare;
databusin[72] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[72] = dontcare;

iaddrbusout[73] = 32'b00000000000000000000001100011000;
instrbusin[73]={ADDI, 5'b00000, 5'b10100, 16'h5544};
daddrbusout[73] = dontcare;
databusin[73] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[73] = dontcare;

iaddrbusout[74] = 32'b00000000000000000000001100011100;
instrbusin[74]={SUBI, 5'b00000, 5'b10100, 16'h5544};
daddrbusout[74] = dontcare;
databusin[74] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[74] = dontcare;

iaddrbusout[75] = 32'b00000000000000000000001100100000;
instrbusin[75]={ADD, 5'b10100, 5'b10100, 5'b10100};
daddrbusout[75] = dontcare;
databusin[75] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[75] = dontcare;

iaddrbusout[76] = 32'b00000000000000000000001100100100;
instrbusin[76]={SLE, 5'b10100, 5'b10100, 5'b10101};
daddrbusout[76] = dontcare;
databusin[76] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[76] = dontcare;

iaddrbusout[77] = 32'b00000000000000000000001100101000;
instrbusin[77]={SLT, 5'b10100, 5'b10100, 5'b10110};
daddrbusout[77] = dontcare;
databusin[77] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[77] = dontcare;

iaddrbusout[78] = 32'b00000000000000000000001100101100;
instrbusin[78]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[78] = dontcare;
databusin[78] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[78] = dontcare;

iaddrbusout[79] = 32'b00000000000000000000001100110000;
instrbusin[79]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[79] = dontcare;
databusin[79] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[79] = dontcare;

iaddrbusout[80] = 32'b00000000000000000000001100110100;
instrbusin[80]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[80] = dontcare;
databusin[80] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[80] = dontcare;

iaddrbusout[81] = 32'b00000000000000000000001100111000;
instrbusin[81]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[81] = dontcare;
databusin[81] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[81] = dontcare;

iaddrbusout[82] = 32'b00000000000000000000001100111100;
instrbusin[82]={SUBI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[82] = dontcare;
databusin[82] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[82] = dontcare;

iaddrbusout[83] = 32'b00000000000000000000001101000000;
instrbusin[83]={SUBI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[83] = dontcare;
databusin[83] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[83] = dontcare;

iaddrbusout[84] = 32'b00000000000000000000001101000100;
instrbusin[84]={SUBI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[84] = dontcare;
databusin[84] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[84] = dontcare;

iaddrbusout[85] = 32'b00000000000000000000001101001000;
instrbusin[85]={XORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[85] = dontcare;
databusin[85] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[85] = dontcare;

iaddrbusout[86] = 32'b00000000000000000000001101001100;
instrbusin[86]={XORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[86] = dontcare;
databusin[86] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[86] = dontcare;

iaddrbusout[87] = 32'b00000000000000000000001101010000;
instrbusin[87]={XORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[87] = dontcare;
databusin[87] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[87] = dontcare;

iaddrbusout[88] = 32'b00000000000000000000001101010100;
instrbusin[88]={ORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[88] = dontcare;
databusin[88] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[88] = dontcare;

iaddrbusout[89] = 32'b00000000000000000000001101011000;
instrbusin[89]={ORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[89] = dontcare;
databusin[89] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[89] = dontcare;

iaddrbusout[90] = 32'b00000000000000000000001101011100;
instrbusin[90]={ORI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[90] = dontcare;
databusin[90] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[90] = dontcare;

iaddrbusout[91] = 32'b00000000000000000000001101100000;
instrbusin[91]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[91] = dontcare;
databusin[91] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[91] = dontcare;

iaddrbusout[92] = 32'b00000000000000000000001101100100;
instrbusin[92]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[92] = dontcare;
databusin[92] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[92] = dontcare;

iaddrbusout[93] = 32'b00000000000000000000001101101000;
instrbusin[93]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[93] = dontcare;
databusin[93] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[93] = dontcare;

iaddrbusout[94] = 32'b00000000000000000000001101101100;
instrbusin[94]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[94] = dontcare;
databusin[94] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[94] = dontcare;

iaddrbusout[95] = 32'b00000000000000000000001101110000;
instrbusin[95]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[95] = dontcare;
databusin[95] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[95] = dontcare;

iaddrbusout[96] = 32'b00000000000000000000001101110100;
instrbusin[96]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[96] = dontcare;
databusin[96] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[96] = dontcare;

iaddrbusout[97] = 32'b00000000000000000000001101111000;
instrbusin[97]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[97] = dontcare;
databusin[97] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[97] = dontcare;

iaddrbusout[98] = 32'b00000000000000000000001101111100;
instrbusin[98]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[98] = dontcare;
databusin[98] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[98] = dontcare;

iaddrbusout[99] = 32'b00000000000000000000001110000000;
instrbusin[99]={ADDI, 5'b00000, 5'b10100, 16'h4444};
daddrbusout[99] = dontcare;
databusin[99] = 32'bzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzzz;
databusout[99] = dontcare;
  
  
// (no. instructions) + (no. loads) + 2*(no. stores) = 35 + 2 + 2*7 = 51
  // 99 + 4 + 2*14 = 131
ntests = 131;
$timeformat(-9,1,"ns",12);
end
//assumes positive edge FF.
//testbench reads databus when clk high, writes databus when clk low.
assign databus = clkd ? 32'bz : databusk;
//Change inputs in middle of period (falling edge).
initial begin
error = 0;
clkd =1;
clk=1;
$display ("Time=%t\n clk=%b", $realtime, clk);
databusk = 32'bz;
//extended reset to set up PC MUX
reset = 1;
$display ("reset=%b", reset);
#5
clk=0;
clkd=0;
$display ("Time=%t\n clk=%b", $realtime, clk);
#5
clk=1;
clkd=1;
$display ("Time=%t\n clk=%b", $realtime, clk);
#5
clk=0;
clkd=0;
$display ("Time=%t\n clk=%b", $realtime, clk);
#5
$display ("Time=%t\n clk=%b", $realtime, clk);
  for (k=0; k<= 99; k=k+1) begin
clk=1;
$display ("Time=%t\n clk=%b", $realtime, clk);
#2
clkd=1;
#3
$display ("Time=%t\n clk=%b", $realtime, clk);
reset = 0;
$display ("reset=%b", reset);
//set load data for 3rd previous instruction
if (k >=3)
databusk = databusin[k-3];
//check PC for this instruction
if (k >= 0) begin
$display (" Testing PC for instruction %d", k);
$display (" Your iaddrbus = %b", iaddrbus);
$display (" Correct iaddrbus = %b", iaddrbusout[k]);
if (iaddrbusout[k] !== iaddrbus) begin
$display (" -------------ERROR. A Mismatch Has Occured-----------");
error = error + 1;
end
end
//put next instruction on ibus
instrbus=instrbusin[k];
$display (" instrbus=%b %b %b %b %b for instruction %d: %s", instrbus[31:26],
instrbus[25:21], instrbus[20:16], instrbus[15:11], instrbus[10:0], k, iname[k]);
//check data address from 3rd previous instruction
if ( (k >= 3) && (daddrbusout[k-3] !== dontcare) ) begin
$display (" Testing data address for instruction %d:", k-3);
$display (" %s", iname[k-3]);
$display (" Your daddrbus = %b", daddrbus);
$display (" Correct daddrbus = %b", daddrbusout[k-3]);
if (daddrbusout[k-3] !== daddrbus) begin
$display (" -------------ERROR. A Mismatch Has Occured-----------");
error = error + 1;
end
end
//check store data from 3rd previous instruction
if ( (k >= 3) && (databusout[k-3] !== dontcare) ) begin
$display (" Testing store data for instruction %d:", k-3);
$display (" %s", iname[k-3]);
$display (" Your databus = %b", databus);
$display (" Correct databus = %b", databusout[k-3]);
if (databusout[k-3] !== databus) begin
$display (" -------------ERROR. A Mismatch Has Occured-----------");
error = error + 1;
end
end
clk = 0;
$display ("Time=%t\n clk=%b", $realtime, clk);
#2
clkd = 0;
#3
$display ("Time=%t\n clk=%b", $realtime, clk);
end
if ( error !== 0) begin
$display("--------- SIMULATION UNSUCCESFUL - MISMATCHES HAVE OCCURED----------");
$display(" No. Of Errors = %d", error);
end
if ( error == 0)
$display("---------YOU DID IT!! SIMULATION SUCCESFULLY FINISHED----------");
end
endmodule
